module config (
	input osc,
);


endmodule